module WB #(parameter WIDTH = 32) (
    input clk,
);



endmodule

